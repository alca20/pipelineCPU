module reg31(data);
	output logic [63:0] data;
	assign data = 0;
endmodule